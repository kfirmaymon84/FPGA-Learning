----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/11/2019 08:17:47 AM
-- Design Name: 
-- Module Name: counter - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use IEEE.std_logic_unsigned.all;
-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity demo_counter is
    Port ( clock : in STD_LOGIC;
           reset : in STD_LOGIC;
           ce : in STD_LOGIC;
           counter : out STD_LOGIC_VECTOR (9 downto 0));
end demo_counter;

architecture Behavioral of demo_counter is
signal count : STD_LOGIC_VECTOR (9 downto 0) := (others => '0');
begin

process (clock)
begin
   if clock='1' and clock'event then
      if reset = '1' then
         count <= (others => '0');
      elsif ce ='1' then
         count <= count + 1;
      end if;
   end if;
end process;

counter <= count;

end Behavioral;
